//// Multiply and Multiply-Add module.

module F_mult (input logic [22:0] a, b 


/// 		MULT MODULE
/// 		46-bit output
/// 	+ nothing	+ Adder
///         |              47-bit out
///         |			|
///	      >ROUNDING UNIT <
