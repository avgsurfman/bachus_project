//// Float mantisa calculator block. Basically a wrapper for other modules. might delete

module 
