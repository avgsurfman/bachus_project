// Priority encoder.

module F_priority_encoder(input logic [22:0] a,
                          output logic [4:0] y);
    always_comb begin
        casez(a)
        23'b00000_0000_0000_0000_0000_00: y=5'd0;
        23'b00000_0000_0000_0000_0000_01: y=5'd1;
        23'b00000_0000_0000_0000_0000_1?: y=5'd2;
        23'b00000_0000_0000_0000_0001_??: y=5'd3;
        23'b00000_0000_0000_0000_001?_??: y=5'd4;
        23'b00000_0000_0000_0000_01??_??: y=5'd5;
        23'b00000_0000_0000_0000_1???_??: y=5'd6;
        23'b00000_0000_0000_0001_????_??: y=5'd7;
        23'b00000_0000_0000_001?_????_??: y=5'd8;
        23'b00000_0000_0000_01??_????_??: y=5'd9;
        23'b00000_0000_0000_1???_????_??: y=5'd10;
        23'b00000_0000_0001_????_????_??: y=5'd11;
        23'b00000_0000_001?_????_????_??: y=5'd12;
        23'b00000_0000_01??_????_????_??: y=5'd13;
        23'b00000_0000_1???_????_????_??: y=5'd14;
        23'b00000_0001_????_????_????_??: y=5'd15;
        23'b00000_001?_????_????_????_??: y=5'd16;
        23'b00000_01??_????_????_????_??: y=5'd17;
        23'b00000_1???_????_????_????_??: y=5'd18;
        23'b00001_????_????_????_????_??: y=5'd19;
        23'b0001?_????_????_????_????_??: y=5'd20;
        23'b001??_????_????_????_????_??: y=5'd21;
        23'b01???_????_????_????_????_??: y=5'd22;
        23'b1????_????_????_????_????_??: y=5'd23;
        endcase
    end
endmodule

