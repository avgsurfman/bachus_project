//// Division Ruine
/// Divider module stub.
module F_div  (input logic [31:0] a, b,
               input logic [2:0]  rounding,  
               //input logic clk,
               output logic flags [4:0], // NV DZ OF UF NX
               output logic [31:0] y);

/// Signal decoders

//// EXP DIFFERENCE


//// MANTISSA division
/// Newton---Raphson goes HERE
// unfortunately this needs batshit fast CSA


//// Exception handling 
/// (can be copied from the mult module)

endmodule
