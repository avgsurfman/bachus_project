//// Multiply module. 
/// TODO: replace with comppressors, specialized prefix adder,
// Fine-tuned 


module F_mult (input logic [22:0] a, b,
              output logic [45:0] mul,
              output logic [4:0] shift_due); 

/// Shift-due uses a priority encoder with casez

endmodule
