//// Division Ruine

module F_div
///     Divider (a, b)
//      Doesn't care about illegal values, just does the computation.
endmodule
