module F_expDiff(input logic [7:0] a, b,
                 output logic [8:0] y);

endmodule
