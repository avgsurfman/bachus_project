//// Top-level file for the FPU.


