//// Add-substract module. 

module F_add (input logic [22:0] a, b 


/// 		ADD MODULE
/// 		24-bit output, sklansky addder
///           Is Special?        
///         Y/return NAN     N/return res
///	      >ROUNDING UNIT <
