//// FPU Regfile.
/// Constains 32 float registers + Float Control-State Register (FCSR).

/// module F_regfile
